`timescale 1ns / 1ps

`define IDX64(x)            ((x) << 6)+:64

// Testbench for the Skein block process implementation
module Skein1024Block_tb;
	
	localparam STARTING_WORK = 2'b00, MIDDLE_SECTION = 2'b01, WAITING_ON_RESULTS = 2'b10;
	genvar x;
	
	// Reg
	reg clk = 1'b0, DataValid = 1'b0;
	
	// Inputs
	reg [1023:0] TestInput;
	reg [1087:0] TestKey;
	reg [191:0] TestType;
	
	always #1 clk = ~clk;
	wire [1023:0] Output;
	wire CompletedSig;
			
    initial
	begin
	
		$dumpfile("SimOutput.lxt2");
		$dumpvars(0, Skein1024Block_tb);
		
		#2;
		
        // Initialize input
        TestInput <= 1024'hA6D8A0A61291CD34F4546149C74CC22E2649339EB37B6519AED442CA29B94FB21BFFD5B90DE16C135743D3A68ED874A160F27B8D098A828BF98FACDB647C0355371E5F0A3B9E81B7F7F78C1BAD4B1DF441B07D5909BE1F3FA16C4845892B8E46A34B94CDB69DFAF73D6E858FC504E56DFD6B3533D9D8B3B11BCECBB3A446FA31;
        TestKey <= 1088'h11409CDB9691AEBB5663952F715D1DDD53D6E4F52E19A6D1FC46DE35C4E2A0860D339D5DAADEE3DC9828030DA0A6388CCC1A9CAFA494DBD30914A20D3DFEA9E49D2599730EF7AB6BB2F6675FA17F0FD23304ACFCA83009983FDBFB11D4A46A3E583A8BFCCE34EB6C6C23C39667038BCAFFCBFE9CA1A2CE265F6E8B1A72F001CA5A4352BE62092156;
        TestType <= 192'h700000000000008070000000000000000000000000000080;

        #2

        // Hold the valid data signal high for one clock cycle
		DataValid <= 1'b1;

		#2;

		DataValid <= 1'b0;

		#2
		
        while(~CompletedSig) #2;
        
        if(Output == 1024'h9078411822E49AAE5512449E8F4ED59107B079C9DF2BCE3971614DDE843E901CBE4AD1BA2E0A2BA8FA2961C972F775C5C6B995F0D482AC8854FC2D17112F99D406C04D28B82118E3852A1A7B236C6C36A6492DF609BD61FC0D6FD0C2F85CB45CD52EBE0DD72D398BFF9AEE231C289271817284E6DBCA4063D96FCEBB0D5AF404)
			$display("PASS.");
		else
			$display("FAIL. 0x%h", Output);

		$finish;
	end
	
	Skein1024Block BlockProcessTest(Output, CompletedSig, clk, DataValid, TestInput, TestKey, TestType);
endmodule
