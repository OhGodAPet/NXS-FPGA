`timescale 1ns / 1ps

`define IDX64(x)            ((x) << 6)+:64

// Testbench for the Skein key injection implementation
// Key is not to be rotated by the injection module
// The round number used is 5.
module SkeinInjectKey_tb;
	
	localparam STARTING_WORK = 2'b00, MIDDLE_SECTION = 2'b01, WAITING_ON_RESULTS = 2'b10;
	genvar x;
	
	// Reg
	reg clk = 1'b0;
	
	// Inputs
	reg [1023:0] TestInput;
	reg [1087:0] TestKey;
	reg [191:0] TestType;
		    
	always #1 clk = ~clk;
	wire [1023:0] Output;
			
    initial
	begin
	
		$dumpfile("SimOutput.lxt2");
		$dumpvars(0, SkeinInjectKey_tb);
		
		#2;
		
        // Initialize input
        TestInput <= 1024'hA6D8A0A61291CD34F4546149C74CC22E2649339EB37B6519AED442CA29B94FB21BFFD5B90DE16C135743D3A68ED874A160F27B8D098A828BF98FACDB647C0355371E5F0A3B9E81B7F7F78C1BAD4B1DF441B07D5909BE1F3FA16C4845892B8E46A34B94CDB69DFAF73D6E858FC504E56DFD6B3533D9D8B3B11BCECBB3A446FA31;
        TestKey <= 1088'h5140285EA2E386F7167680BE7897F81971A3086ACC6CC8F057C1D69EA96127F3ABB56DF877FDECB8B1E9D263648DBE76F3CB2FA1739B5285E2AB244823C589F99B9F238E28F0C967101D5D42065C65273E274D718830E81ED86F7A18605FB3D75E674880CB9E47A4797A1003D479B77B3E245EDF8787BF9EAB986FFFA8FEF30A34646120A8B4C7D4;
        TestType <= 192'hCD4818BC80D049A3AA3F44C0CBE08F9C242E7683A3E1B23C;
        #2;
        #2;

        if(Output == 1024'hA6D8A0A61291CD391882D7CD6B2E746AF3914C5B344BAEBC5A89B0C2A1B73C6ACDE9A81C726F2A894B0F03480273C726439D9FD52D500C84952ED0698D6CCCBC473BBC4C41FAE6DE361ED98D357C06121A1FF7716A1DD316FFD390C654C9D5EA1CC5A4D18B17B2727B92E46F4C8CA50BA903A53382D7A6BB50332CD44CFBC205)
			$display("PASS.");
		else
			$display("FAIL. 0x%h", Output);

		$finish;
	end
	
	SkeinInjectKey #(.RNDNUM(5), .RNDNUM_MOD_3(2)) TestInjection(Output, clk, TestInput, TestKey, TestType);
endmodule
